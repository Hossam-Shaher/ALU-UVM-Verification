`ifndef ALU_SEQUENCER_SV
  `define ALU_SEQUENCER_SV

  typedef class alu_seq_item_drv;

  typedef uvm_sequencer#(alu_seq_item_drv) alu_sequencer; 

`endif //ALU_SEQUENCER_SV